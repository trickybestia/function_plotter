`timescale 1ns / 1ps

module stack_machine_tb;

reg clk;
   
endmodule
