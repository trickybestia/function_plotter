`timescale 1ns / 1ps

module parser_tb;

reg clk;
   
endmodule
